`timescale 1ns/1ps
module DSP48A1_tb();

